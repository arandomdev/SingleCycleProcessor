`timescale 1ns / 1ns

package TopTestVectors;
  typedef struct {
    string  name;
    string  instructionsFile;
    integer initialRegFileState[31];  // Excludes x0
    integer finalRegFileState[31];    // Excludes x0
    integer initialRamState[256];
    integer finalRamState[256];
  } test_vector_t;

  test_vector_t testVectors[] = '{
      '{
          name: "Program 1",
          instructionsFile: "program1.mem",
          initialRegFileState: '{31{32'h00000000}},
          finalRegFileState: '{
              32'h00000000,
              32'h00000010,
              32'h00000064,
              32'h00000008,
              32'h00000010,
              32'h0000006c,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          initialRamState: '{256{32'h00000000}},
          finalRamState: '{
              32'h00000010,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h0000006c,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          }
      },
      '{
          name: "Program 2",
          instructionsFile: "program2.mem",
          initialRegFileState: '{31{32'h00000000}},
          finalRegFileState: '{
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h0000000c,
              32'h0000000f,
              32'h00000017,
              32'h00000000,
              32'h000000a1,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000248,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000007,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          initialRamState: '{256{32'h00000000}},
          finalRamState: '{
              32'h00000000,
              32'h00000000,
              32'h0000000f,
              32'h00000248,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          }
      },
      '{
          name: "Program 3",
          instructionsFile: "program3.mem",
          initialRegFileState: '{
              32'h00000000,
              32'h000000fc,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          finalRegFileState: '{
              32'h00000008,
              32'h000000fc,
              32'h00000000,
              32'h00000000,
              32'h02611500,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h1c8cfc00,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          initialRamState: '{256{32'h00000000}},
          finalRamState: '{
              32'h1c8cfc00,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000001,
              32'h00000034,
              32'h00000002,
              32'h00000034,
              32'h00000003,
              32'h00000034,
              32'h00000004,
              32'h00000034,
              32'h00000005,
              32'h00000034,
              32'h00000006,
              32'h00000034,
              32'h00000007,
              32'h00000034,
              32'h00000008,
              32'h00000034,
              32'h00000009,
              32'h00000034,
              32'h0000000a,
              32'h00000034,
              32'h0000000b,
              32'h00000034,
              32'h0000000c,
              32'h00000008,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          }
      },
      '{
          name: "Program 4",
          instructionsFile: "program4.mem",
          initialRegFileState: '{31{32'h00000000}},
          finalRegFileState: '{
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000015,
              32'h00000007,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000005,
              32'h00000018,
              32'h00000005,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          initialRamState: '{
              32'h00000005,
              32'h00000002,
              32'h00000006,
              32'h00000005,
              32'h00000001,
              32'h00000007,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          finalRamState: '{
              32'h00000005,
              32'h00000002,
              32'h00000006,
              32'h00000005,
              32'h00000001,
              32'h00000007,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          }
      }
  };
endpackage
