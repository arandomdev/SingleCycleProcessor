`timescale 1ns / 1ns

package TopTestVectors;
  typedef struct {
    string name;
    int instructions[];
    integer initialRegFileState[31];  // Excludes x0
    integer finalRegFileState[31];  // Excludes x0
    integer initialRamState[256];
    integer finalRamState[256];
  } test_vector_t;

  test_vector_t testVectors[] = '{
      '{
          name: "Program 1",
          instructions: '{
              32'h00000093,  // addi x1, x0, 0
              32'h01000113,  // addi x2, x0, 16
              32'h06400193,  // addi x3, x0, 100
              32'h00800213,  // addi x4, x0, 8
              32'h002082b3,  // add x5, x1, x2
              32'h00418333,  // add x6, x3, x4
              32'h0050a023,  // sw x5, 0(x1)
              32'h00612223,  // sw x6, 4(x2)
              32'h0000007f  // HALT
          },
          initialRegFileState: '{31{32'h00000000}},
          finalRegFileState: '{
              32'h00000000,
              32'h00000010,
              32'h00000064,
              32'h00000008,
              32'h00000010,
              32'h0000006c,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          initialRamState: '{256{32'h00000000}},
          finalRamState: '{
              32'h00000010,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h0000006c,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          }
      },
      '{
          name: "Program 2",
          instructions: '{
              32'h00800293,  // addi t0, x0, 8
              32'h00f00313,  // addi t1, x0, 15
              32'h0062a023,  // sw t1, 0(t0)
              32'h005303b3,  // add t2, t1, t0
              32'h40530e33,  // sub t3, t1, t0
              32'h03c384b3,  // mul s1, t2, t3
              32'h00428293,  // addi t0, t0, 4
              32'hffc2a903,  // lw s2, -4(t0)
              32'h41248933,  // sub s2, s1, s2
              32'h00291913,  // slli s2, s2, 2
              32'h0122a023,  // sw s2, 0(t0)
              32'h0000007f  // HALT
          },
          initialRegFileState: '{31{32'h00000000}},
          finalRegFileState: '{
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h0000000c,
              32'h0000000f,
              32'h00000017,
              32'h00000000,
              32'h000000a1,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000248,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000007,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          initialRamState: '{256{32'h00000000}},
          finalRamState: '{
              32'h00000000,
              32'h00000000,
              32'h0000000f,
              32'h00000248,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          }
      },
      '{
          name: "Program 3",
          instructions: '{
              32'h00c00513,  // addi a0, x0, 12
              32'h00c000ef,  // jal ra, fact
              32'h00a02023,  // sw a0, 0(x0)
              32'h0000007f,  // HALT
              32'hff810113,  // fact: addi sp, sp, -8
              32'h00112223,  // sw ra, 4(sp)
              32'h00a12023,  // sw a0, 0(sp)
              32'hfff50513,  // addi a0, a0, -1
              32'h00051863,  // bne a0, x0, else
              32'h00100513,  // addi a0, x0, 1
              32'h00810113,  // addi sp, sp, 8
              32'h00008067,  // jalr x0, 0(ra)
              32'hfe1ff0ef,  // else: jal ra, fact
              32'h00050293,  // addi t0, a0,0
              32'h00012503,  // lw a0, 0(sp)
              32'h00412083,  // lw ra, 4(sp)
              32'h00810113,  // addi sp, sp, 8
              32'h02550533,  // mul a0, a0, t0
              32'h00008067  // jalr x0, 0(ra)
          },
          initialRegFileState: '{
              32'h00000000,
              32'h000000fc,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          finalRegFileState: '{
              32'h00000008,
              32'h000000fc,
              32'h00000000,
              32'h00000000,
              32'h02611500,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h1c8cfc00,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          },
          initialRamState: '{256{32'h00000000}},
          finalRamState: '{
              32'h1c8cfc00,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000001,
              32'h00000034,
              32'h00000002,
              32'h00000034,
              32'h00000003,
              32'h00000034,
              32'h00000004,
              32'h00000034,
              32'h00000005,
              32'h00000034,
              32'h00000006,
              32'h00000034,
              32'h00000007,
              32'h00000034,
              32'h00000008,
              32'h00000034,
              32'h00000009,
              32'h00000034,
              32'h0000000a,
              32'h00000034,
              32'h0000000b,
              32'h00000034,
              32'h0000000c,
              32'h00000008,
              32'h00000000,
              32'h00000000,
              32'h00000000,
              32'h00000000
          }
      }
  };
endpackage
